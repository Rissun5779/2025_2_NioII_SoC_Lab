
module Nios2 (
	clk_clk,
	reset_reset_n,
	pio_led_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[9:0]	pio_led_export;
endmodule
