
module Nios2 (
	clk_clk,
	pio_led_export,
	reset_reset_n);	

	input		clk_clk;
	output	[9:0]	pio_led_export;
	input		reset_reset_n;
endmodule
