-- nios2.vhd

-- Generated using ACDS version 13.1 162 at 2026.02.27.22:37:12

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2 is
	port (
		clk_clk        : in  std_logic                    := '0'; --     clk.clk
		led_pio_export : out std_logic_vector(7 downto 0);        -- led_pio.export
		reset_reset_n  : in  std_logic                    := '0'  --   reset.reset_n
	);
end entity nios2;

architecture rtl of nios2 is
	component nios2_nios2 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(17 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios2_nios2;

	component nios2_RAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios2_RAM;

	component nios2_JUART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios2_JUART;

	component nios2_LED_PIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios2_LED_PIO;

	component nios2_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			nios2_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_data_master_address                 : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			JUART_avalon_jtag_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			JUART_avalon_jtag_slave_write             : out std_logic;                                        -- write
			JUART_avalon_jtag_slave_read              : out std_logic;                                        -- read
			JUART_avalon_jtag_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JUART_avalon_jtag_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			JUART_avalon_jtag_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			JUART_avalon_jtag_slave_chipselect        : out std_logic;                                        -- chipselect
			LED_PIO_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			LED_PIO_s1_write                          : out std_logic;                                        -- write
			LED_PIO_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LED_PIO_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			LED_PIO_s1_chipselect                     : out std_logic;                                        -- chipselect
			nios2_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			RAM_s1_address                            : out std_logic_vector(13 downto 0);                    -- address
			RAM_s1_write                              : out std_logic;                                        -- write
			RAM_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			RAM_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM_s1_chipselect                         : out std_logic;                                        -- chipselect
			RAM_s1_clken                              : out std_logic                                         -- clken
		);
	end component nios2_mm_interconnect_0;

	component nios2_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal mm_interconnect_0_led_pio_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:LED_PIO_s1_writedata -> LED_PIO:writedata
	signal mm_interconnect_0_led_pio_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LED_PIO_s1_address -> LED_PIO:address
	signal mm_interconnect_0_led_pio_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:LED_PIO_s1_chipselect -> LED_PIO:chipselect
	signal mm_interconnect_0_led_pio_s1_write                        : std_logic;                     -- mm_interconnect_0:LED_PIO_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_readdata                     : std_logic_vector(31 downto 0); -- LED_PIO:readdata -> mm_interconnect_0:LED_PIO_s1_readdata
	signal mm_interconnect_0_juart_avalon_jtag_slave_waitrequest     : std_logic;                     -- JUART:av_waitrequest -> mm_interconnect_0:JUART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_juart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JUART_avalon_jtag_slave_writedata -> JUART:av_writedata
	signal mm_interconnect_0_juart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JUART_avalon_jtag_slave_address -> JUART:av_address
	signal mm_interconnect_0_juart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JUART_avalon_jtag_slave_chipselect -> JUART:av_chipselect
	signal mm_interconnect_0_juart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JUART_avalon_jtag_slave_write -> mm_interconnect_0_juart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_juart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JUART_avalon_jtag_slave_read -> mm_interconnect_0_juart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_juart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JUART:av_readdata -> mm_interconnect_0:JUART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_nios2_jtag_debug_module_waitrequest     : std_logic;                     -- nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_jtag_debug_module_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	signal mm_interconnect_0_nios2_jtag_debug_module_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	signal mm_interconnect_0_nios2_jtag_debug_module_write           : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	signal mm_interconnect_0_nios2_jtag_debug_module_read            : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	signal mm_interconnect_0_nios2_jtag_debug_module_readdata        : std_logic_vector(31 downto 0); -- nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_jtag_debug_module_debugaccess     : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_jtag_debug_module_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	signal nios2_data_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_writedata                               : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	signal nios2_data_master_address                                 : std_logic_vector(17 downto 0); -- nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	signal nios2_data_master_write                                   : std_logic;                     -- nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	signal nios2_data_master_read                                    : std_logic;                     -- nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	signal nios2_data_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_debugaccess                             : std_logic;                     -- nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	signal nios2_data_master_byteenable                              : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	signal mm_interconnect_0_ram_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	signal mm_interconnect_0_ram_s1_address                          : std_logic_vector(13 downto 0); -- mm_interconnect_0:RAM_s1_address -> RAM:address
	signal mm_interconnect_0_ram_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	signal mm_interconnect_0_ram_s1_clken                            : std_logic;                     -- mm_interconnect_0:RAM_s1_clken -> RAM:clken
	signal mm_interconnect_0_ram_s1_write                            : std_logic;                     -- mm_interconnect_0:RAM_s1_write -> RAM:write
	signal mm_interconnect_0_ram_s1_readdata                         : std_logic_vector(31 downto 0); -- RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	signal mm_interconnect_0_ram_s1_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	signal nios2_instruction_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                          : std_logic_vector(17 downto 0); -- nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	signal nios2_instruction_master_read                             : std_logic;                     -- nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	signal nios2_instruction_master_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	signal irq_mapper_receiver0_irq                                  : std_logic;                     -- JUART:av_irq -> irq_mapper:receiver0_irq
	signal nios2_d_irq_irq                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:d_irq
	signal rst_controller_reset_out_reset                            : std_logic;                     -- rst_controller:reset_out -> [RAM:reset, irq_mapper:reset, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                        : std_logic;                     -- rst_controller:reset_req -> [RAM:reset_req, nios2:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                   : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_led_pio_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> LED_PIO:write_n
	signal mm_interconnect_0_juart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_juart_avalon_jtag_slave_write:inv -> JUART:av_write_n
	signal mm_interconnect_0_juart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_juart_avalon_jtag_slave_read:inv -> JUART:av_read_n
	signal rst_controller_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JUART:rst_n, LED_PIO:reset_n, nios2:reset_n]

begin

	nios2 : component nios2_nios2
		port map (
			clk                                   => clk_clk,                                               --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,              --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                             => nios2_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_data_master_read,                                --                          .read
			d_readdata                            => nios2_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_data_master_write,                               --                          .write
			d_writedata                           => nios2_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                  --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                   -- custom_instruction_master.readra
		);

	ram : component nios2_RAM
		port map (
			clk        => clk_clk,                             --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req   --       .reset_req
		);

	juart : component nios2_JUART
		port map (
			clk            => clk_clk,                                                   --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_juart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_juart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_juart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_juart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_juart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_juart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_juart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                   --               irq.irq
		);

	led_pio : component nios2_LED_PIO
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_export                                -- external_connection.export
		);

	mm_interconnect_0 : component nios2_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                               --                           clk_0_clk.clk
			nios2_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                        -- nios2_reset_n_reset_bridge_in_reset.reset
			nios2_data_master_address                 => nios2_data_master_address,                             --                   nios2_data_master.address
			nios2_data_master_waitrequest             => nios2_data_master_waitrequest,                         --                                    .waitrequest
			nios2_data_master_byteenable              => nios2_data_master_byteenable,                          --                                    .byteenable
			nios2_data_master_read                    => nios2_data_master_read,                                --                                    .read
			nios2_data_master_readdata                => nios2_data_master_readdata,                            --                                    .readdata
			nios2_data_master_write                   => nios2_data_master_write,                               --                                    .write
			nios2_data_master_writedata               => nios2_data_master_writedata,                           --                                    .writedata
			nios2_data_master_debugaccess             => nios2_data_master_debugaccess,                         --                                    .debugaccess
			nios2_instruction_master_address          => nios2_instruction_master_address,                      --            nios2_instruction_master.address
			nios2_instruction_master_waitrequest      => nios2_instruction_master_waitrequest,                  --                                    .waitrequest
			nios2_instruction_master_read             => nios2_instruction_master_read,                         --                                    .read
			nios2_instruction_master_readdata         => nios2_instruction_master_readdata,                     --                                    .readdata
			JUART_avalon_jtag_slave_address           => mm_interconnect_0_juart_avalon_jtag_slave_address,     --             JUART_avalon_jtag_slave.address
			JUART_avalon_jtag_slave_write             => mm_interconnect_0_juart_avalon_jtag_slave_write,       --                                    .write
			JUART_avalon_jtag_slave_read              => mm_interconnect_0_juart_avalon_jtag_slave_read,        --                                    .read
			JUART_avalon_jtag_slave_readdata          => mm_interconnect_0_juart_avalon_jtag_slave_readdata,    --                                    .readdata
			JUART_avalon_jtag_slave_writedata         => mm_interconnect_0_juart_avalon_jtag_slave_writedata,   --                                    .writedata
			JUART_avalon_jtag_slave_waitrequest       => mm_interconnect_0_juart_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			JUART_avalon_jtag_slave_chipselect        => mm_interconnect_0_juart_avalon_jtag_slave_chipselect,  --                                    .chipselect
			LED_PIO_s1_address                        => mm_interconnect_0_led_pio_s1_address,                  --                          LED_PIO_s1.address
			LED_PIO_s1_write                          => mm_interconnect_0_led_pio_s1_write,                    --                                    .write
			LED_PIO_s1_readdata                       => mm_interconnect_0_led_pio_s1_readdata,                 --                                    .readdata
			LED_PIO_s1_writedata                      => mm_interconnect_0_led_pio_s1_writedata,                --                                    .writedata
			LED_PIO_s1_chipselect                     => mm_interconnect_0_led_pio_s1_chipselect,               --                                    .chipselect
			nios2_jtag_debug_module_address           => mm_interconnect_0_nios2_jtag_debug_module_address,     --             nios2_jtag_debug_module.address
			nios2_jtag_debug_module_write             => mm_interconnect_0_nios2_jtag_debug_module_write,       --                                    .write
			nios2_jtag_debug_module_read              => mm_interconnect_0_nios2_jtag_debug_module_read,        --                                    .read
			nios2_jtag_debug_module_readdata          => mm_interconnect_0_nios2_jtag_debug_module_readdata,    --                                    .readdata
			nios2_jtag_debug_module_writedata         => mm_interconnect_0_nios2_jtag_debug_module_writedata,   --                                    .writedata
			nios2_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_jtag_debug_module_byteenable,  --                                    .byteenable
			nios2_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_jtag_debug_module_waitrequest, --                                    .waitrequest
			nios2_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_jtag_debug_module_debugaccess, --                                    .debugaccess
			RAM_s1_address                            => mm_interconnect_0_ram_s1_address,                      --                              RAM_s1.address
			RAM_s1_write                              => mm_interconnect_0_ram_s1_write,                        --                                    .write
			RAM_s1_readdata                           => mm_interconnect_0_ram_s1_readdata,                     --                                    .readdata
			RAM_s1_writedata                          => mm_interconnect_0_ram_s1_writedata,                    --                                    .writedata
			RAM_s1_byteenable                         => mm_interconnect_0_ram_s1_byteenable,                   --                                    .byteenable
			RAM_s1_chipselect                         => mm_interconnect_0_ram_s1_chipselect,                   --                                    .chipselect
			RAM_s1_clken                              => mm_interconnect_0_ram_s1_clken                         --                                    .clken
		);

	irq_mapper : component nios2_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_d_irq_irq                 --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_juart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_juart_avalon_jtag_slave_write;

	mm_interconnect_0_juart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_juart_avalon_jtag_slave_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios2
