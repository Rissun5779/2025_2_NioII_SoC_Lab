// nios2.v

// Generated using ACDS version 13.1 162 at 2026.02.27.22:37:49

`timescale 1 ps / 1 ps
module nios2 (
		input  wire       clk_clk,        //     clk.clk
		output wire [7:0] led_pio_export, // led_pio.export
		input  wire       reset_reset_n   //   reset.reset_n
	);

	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                    // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire  [13:0] mm_interconnect_0_ram_s1_address;                      // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire         mm_interconnect_0_ram_s1_chipselect;                   // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire         mm_interconnect_0_ram_s1_clken;                        // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_ram_s1_write;                        // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                     // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                   // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_juart_avalon_jtag_slave_waitrequest; // JUART:av_waitrequest -> mm_interconnect_0:JUART_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_juart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JUART_avalon_jtag_slave_writedata -> JUART:av_writedata
	wire   [0:0] mm_interconnect_0_juart_avalon_jtag_slave_address;     // mm_interconnect_0:JUART_avalon_jtag_slave_address -> JUART:av_address
	wire         mm_interconnect_0_juart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JUART_avalon_jtag_slave_chipselect -> JUART:av_chipselect
	wire         mm_interconnect_0_juart_avalon_jtag_slave_write;       // mm_interconnect_0:JUART_avalon_jtag_slave_write -> JUART:av_write_n
	wire         mm_interconnect_0_juart_avalon_jtag_slave_read;        // mm_interconnect_0:JUART_avalon_jtag_slave_read -> JUART:av_read_n
	wire  [31:0] mm_interconnect_0_juart_avalon_jtag_slave_readdata;    // JUART:av_readdata -> mm_interconnect_0:JUART_avalon_jtag_slave_readdata
	wire         nios2_data_master_waitrequest;                         // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                           // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [17:0] nios2_data_master_address;                             // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                               // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                            // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                         // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire   [3:0] nios2_data_master_byteenable;                          // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [17:0] nios2_instruction_master_address;                      // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                         // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                     // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                // mm_interconnect_0:LED_PIO_s1_writedata -> LED_PIO:writedata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                  // mm_interconnect_0:LED_PIO_s1_address -> LED_PIO:address
	wire         mm_interconnect_0_led_pio_s1_chipselect;               // mm_interconnect_0:LED_PIO_s1_chipselect -> LED_PIO:chipselect
	wire         mm_interconnect_0_led_pio_s1_write;                    // mm_interconnect_0:LED_PIO_s1_write -> LED_PIO:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                 // LED_PIO:readdata -> mm_interconnect_0:LED_PIO_s1_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest; // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;     // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;       // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;        // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;    // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                              // JUART:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [JUART:rst_n, LED_PIO:reset_n, RAM:reset, irq_mapper:reset, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [RAM:reset_req, nios2:reset_req, rst_translator:reset_req_in]

	nios2_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                      //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	nios2_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)   //       .reset_req
	);

	nios2_JUART juart (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_juart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_juart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_juart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_juart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_juart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_juart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_juart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	nios2_LED_PIO led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	nios2_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                               //                           clk_0_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                 (nios2_data_master_address),                             //                   nios2_data_master.address
		.nios2_data_master_waitrequest             (nios2_data_master_waitrequest),                         //                                    .waitrequest
		.nios2_data_master_byteenable              (nios2_data_master_byteenable),                          //                                    .byteenable
		.nios2_data_master_read                    (nios2_data_master_read),                                //                                    .read
		.nios2_data_master_readdata                (nios2_data_master_readdata),                            //                                    .readdata
		.nios2_data_master_write                   (nios2_data_master_write),                               //                                    .write
		.nios2_data_master_writedata               (nios2_data_master_writedata),                           //                                    .writedata
		.nios2_data_master_debugaccess             (nios2_data_master_debugaccess),                         //                                    .debugaccess
		.nios2_instruction_master_address          (nios2_instruction_master_address),                      //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                  //                                    .waitrequest
		.nios2_instruction_master_read             (nios2_instruction_master_read),                         //                                    .read
		.nios2_instruction_master_readdata         (nios2_instruction_master_readdata),                     //                                    .readdata
		.JUART_avalon_jtag_slave_address           (mm_interconnect_0_juart_avalon_jtag_slave_address),     //             JUART_avalon_jtag_slave.address
		.JUART_avalon_jtag_slave_write             (mm_interconnect_0_juart_avalon_jtag_slave_write),       //                                    .write
		.JUART_avalon_jtag_slave_read              (mm_interconnect_0_juart_avalon_jtag_slave_read),        //                                    .read
		.JUART_avalon_jtag_slave_readdata          (mm_interconnect_0_juart_avalon_jtag_slave_readdata),    //                                    .readdata
		.JUART_avalon_jtag_slave_writedata         (mm_interconnect_0_juart_avalon_jtag_slave_writedata),   //                                    .writedata
		.JUART_avalon_jtag_slave_waitrequest       (mm_interconnect_0_juart_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.JUART_avalon_jtag_slave_chipselect        (mm_interconnect_0_juart_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.LED_PIO_s1_address                        (mm_interconnect_0_led_pio_s1_address),                  //                          LED_PIO_s1.address
		.LED_PIO_s1_write                          (mm_interconnect_0_led_pio_s1_write),                    //                                    .write
		.LED_PIO_s1_readdata                       (mm_interconnect_0_led_pio_s1_readdata),                 //                                    .readdata
		.LED_PIO_s1_writedata                      (mm_interconnect_0_led_pio_s1_writedata),                //                                    .writedata
		.LED_PIO_s1_chipselect                     (mm_interconnect_0_led_pio_s1_chipselect),               //                                    .chipselect
		.nios2_jtag_debug_module_address           (mm_interconnect_0_nios2_jtag_debug_module_address),     //             nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write             (mm_interconnect_0_nios2_jtag_debug_module_write),       //                                    .write
		.nios2_jtag_debug_module_read              (mm_interconnect_0_nios2_jtag_debug_module_read),        //                                    .read
		.nios2_jtag_debug_module_readdata          (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                                    .readdata
		.nios2_jtag_debug_module_writedata         (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                                    .writedata
		.nios2_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                                    .byteenable
		.nios2_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                                    .waitrequest
		.nios2_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                                    .debugaccess
		.RAM_s1_address                            (mm_interconnect_0_ram_s1_address),                      //                              RAM_s1.address
		.RAM_s1_write                              (mm_interconnect_0_ram_s1_write),                        //                                    .write
		.RAM_s1_readdata                           (mm_interconnect_0_ram_s1_readdata),                     //                                    .readdata
		.RAM_s1_writedata                          (mm_interconnect_0_ram_s1_writedata),                    //                                    .writedata
		.RAM_s1_byteenable                         (mm_interconnect_0_ram_s1_byteenable),                   //                                    .byteenable
		.RAM_s1_chipselect                         (mm_interconnect_0_ram_s1_chipselect),                   //                                    .chipselect
		.RAM_s1_clken                              (mm_interconnect_0_ram_s1_clken)                         //                                    .clken
	);

	nios2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
